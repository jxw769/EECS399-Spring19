// test1a.v

// Generated using ACDS version 17.0 595

`timescale 1 ps / 1 ps
module test1a (
		output wire [7:0]  addr_external_connection_export,       //       addr_external_connection.export
		input  wire        clk_clk,                               //                            clk.clk
		input  wire        done_external_connection_export,       //       done_external_connection.export
		output wire [7:0]  gpio_external_connection_export,       //       gpio_external_connection.export
		output wire [7:0]  led_external_connection_export,        //        led_external_connection.export
		output wire        m_reset_external_connection_export,    //    m_reset_external_connection.export
		output wire        oper_external_connection_export,       //       oper_external_connection.export
		input  wire        reset_reset_n,                         //                          reset.reset_n
		output wire        start_16_external_connection_export,   //   start_16_external_connection.export
		output wire        start_external_connection_export,      //      start_external_connection.export
		output wire [15:0] wr_data_16_external_connection_export, // wr_data_16_external_connection.export
		output wire [31:0] wr_data_external_connection_export     //    wr_data_external_connection.export
	);

	wire  [31:0] master_0_master_readdata;                   // mm_interconnect_0:master_0_master_readdata -> master_0:master_readdata
	wire         master_0_master_waitrequest;                // mm_interconnect_0:master_0_master_waitrequest -> master_0:master_waitrequest
	wire  [31:0] master_0_master_address;                    // master_0:master_address -> mm_interconnect_0:master_0_master_address
	wire         master_0_master_read;                       // master_0:master_read -> mm_interconnect_0:master_0_master_read
	wire   [3:0] master_0_master_byteenable;                 // master_0:master_byteenable -> mm_interconnect_0:master_0_master_byteenable
	wire         master_0_master_readdatavalid;              // mm_interconnect_0:master_0_master_readdatavalid -> master_0:master_readdatavalid
	wire         master_0_master_write;                      // master_0:master_write -> mm_interconnect_0:master_0_master_write
	wire  [31:0] master_0_master_writedata;                  // master_0:master_writedata -> mm_interconnect_0:master_0_master_writedata
	wire         mm_interconnect_0_led_s1_chipselect;        // mm_interconnect_0:LED_s1_chipselect -> LED:chipselect
	wire  [31:0] mm_interconnect_0_led_s1_readdata;          // LED:readdata -> mm_interconnect_0:LED_s1_readdata
	wire   [1:0] mm_interconnect_0_led_s1_address;           // mm_interconnect_0:LED_s1_address -> LED:address
	wire         mm_interconnect_0_led_s1_write;             // mm_interconnect_0:LED_s1_write -> LED:write_n
	wire  [31:0] mm_interconnect_0_led_s1_writedata;         // mm_interconnect_0:LED_s1_writedata -> LED:writedata
	wire         mm_interconnect_0_addr_s1_chipselect;       // mm_interconnect_0:ADDR_s1_chipselect -> ADDR:chipselect
	wire  [31:0] mm_interconnect_0_addr_s1_readdata;         // ADDR:readdata -> mm_interconnect_0:ADDR_s1_readdata
	wire   [1:0] mm_interconnect_0_addr_s1_address;          // mm_interconnect_0:ADDR_s1_address -> ADDR:address
	wire         mm_interconnect_0_addr_s1_write;            // mm_interconnect_0:ADDR_s1_write -> ADDR:write_n
	wire  [31:0] mm_interconnect_0_addr_s1_writedata;        // mm_interconnect_0:ADDR_s1_writedata -> ADDR:writedata
	wire         mm_interconnect_0_wr_data_s1_chipselect;    // mm_interconnect_0:WR_DATA_s1_chipselect -> WR_DATA:chipselect
	wire  [31:0] mm_interconnect_0_wr_data_s1_readdata;      // WR_DATA:readdata -> mm_interconnect_0:WR_DATA_s1_readdata
	wire   [1:0] mm_interconnect_0_wr_data_s1_address;       // mm_interconnect_0:WR_DATA_s1_address -> WR_DATA:address
	wire         mm_interconnect_0_wr_data_s1_write;         // mm_interconnect_0:WR_DATA_s1_write -> WR_DATA:write_n
	wire  [31:0] mm_interconnect_0_wr_data_s1_writedata;     // mm_interconnect_0:WR_DATA_s1_writedata -> WR_DATA:writedata
	wire         mm_interconnect_0_gpio_s1_chipselect;       // mm_interconnect_0:GPIO_s1_chipselect -> GPIO:chipselect
	wire  [31:0] mm_interconnect_0_gpio_s1_readdata;         // GPIO:readdata -> mm_interconnect_0:GPIO_s1_readdata
	wire   [1:0] mm_interconnect_0_gpio_s1_address;          // mm_interconnect_0:GPIO_s1_address -> GPIO:address
	wire         mm_interconnect_0_gpio_s1_write;            // mm_interconnect_0:GPIO_s1_write -> GPIO:write_n
	wire  [31:0] mm_interconnect_0_gpio_s1_writedata;        // mm_interconnect_0:GPIO_s1_writedata -> GPIO:writedata
	wire         mm_interconnect_0_start_s1_chipselect;      // mm_interconnect_0:START_s1_chipselect -> START:chipselect
	wire  [31:0] mm_interconnect_0_start_s1_readdata;        // START:readdata -> mm_interconnect_0:START_s1_readdata
	wire   [1:0] mm_interconnect_0_start_s1_address;         // mm_interconnect_0:START_s1_address -> START:address
	wire         mm_interconnect_0_start_s1_write;           // mm_interconnect_0:START_s1_write -> START:write_n
	wire  [31:0] mm_interconnect_0_start_s1_writedata;       // mm_interconnect_0:START_s1_writedata -> START:writedata
	wire         mm_interconnect_0_oper_s1_chipselect;       // mm_interconnect_0:OPER_s1_chipselect -> OPER:chipselect
	wire  [31:0] mm_interconnect_0_oper_s1_readdata;         // OPER:readdata -> mm_interconnect_0:OPER_s1_readdata
	wire   [1:0] mm_interconnect_0_oper_s1_address;          // mm_interconnect_0:OPER_s1_address -> OPER:address
	wire         mm_interconnect_0_oper_s1_write;            // mm_interconnect_0:OPER_s1_write -> OPER:write_n
	wire  [31:0] mm_interconnect_0_oper_s1_writedata;        // mm_interconnect_0:OPER_s1_writedata -> OPER:writedata
	wire  [31:0] mm_interconnect_0_done_s1_readdata;         // DONE:readdata -> mm_interconnect_0:DONE_s1_readdata
	wire   [1:0] mm_interconnect_0_done_s1_address;          // mm_interconnect_0:DONE_s1_address -> DONE:address
	wire         mm_interconnect_0_m_reset_s1_chipselect;    // mm_interconnect_0:M_RESET_s1_chipselect -> M_RESET:chipselect
	wire  [31:0] mm_interconnect_0_m_reset_s1_readdata;      // M_RESET:readdata -> mm_interconnect_0:M_RESET_s1_readdata
	wire   [1:0] mm_interconnect_0_m_reset_s1_address;       // mm_interconnect_0:M_RESET_s1_address -> M_RESET:address
	wire         mm_interconnect_0_m_reset_s1_write;         // mm_interconnect_0:M_RESET_s1_write -> M_RESET:write_n
	wire  [31:0] mm_interconnect_0_m_reset_s1_writedata;     // mm_interconnect_0:M_RESET_s1_writedata -> M_RESET:writedata
	wire         mm_interconnect_0_wr_data_16_s1_chipselect; // mm_interconnect_0:WR_DATA_16_s1_chipselect -> WR_DATA_16:chipselect
	wire  [31:0] mm_interconnect_0_wr_data_16_s1_readdata;   // WR_DATA_16:readdata -> mm_interconnect_0:WR_DATA_16_s1_readdata
	wire   [1:0] mm_interconnect_0_wr_data_16_s1_address;    // mm_interconnect_0:WR_DATA_16_s1_address -> WR_DATA_16:address
	wire         mm_interconnect_0_wr_data_16_s1_write;      // mm_interconnect_0:WR_DATA_16_s1_write -> WR_DATA_16:write_n
	wire  [31:0] mm_interconnect_0_wr_data_16_s1_writedata;  // mm_interconnect_0:WR_DATA_16_s1_writedata -> WR_DATA_16:writedata
	wire         mm_interconnect_0_start_16_s1_chipselect;   // mm_interconnect_0:START_16_s1_chipselect -> START_16:chipselect
	wire  [31:0] mm_interconnect_0_start_16_s1_readdata;     // START_16:readdata -> mm_interconnect_0:START_16_s1_readdata
	wire   [1:0] mm_interconnect_0_start_16_s1_address;      // mm_interconnect_0:START_16_s1_address -> START_16:address
	wire         mm_interconnect_0_start_16_s1_write;        // mm_interconnect_0:START_16_s1_write -> START_16:write_n
	wire  [31:0] mm_interconnect_0_start_16_s1_writedata;    // mm_interconnect_0:START_16_s1_writedata -> START_16:writedata
	wire         rst_controller_reset_out_reset;             // rst_controller:reset_out -> [ADDR:reset_n, DONE:reset_n, GPIO:reset_n, LED:reset_n, M_RESET:reset_n, OPER:reset_n, START:reset_n, START_16:reset_n, WR_DATA:reset_n, WR_DATA_16:reset_n, mm_interconnect_0:LED_reset_reset_bridge_in_reset_reset, mm_interconnect_0:master_0_clk_reset_reset_bridge_in_reset_reset]

	test1a_ADDR addr (
		.clk        (clk_clk),                              //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),      //               reset.reset_n
		.address    (mm_interconnect_0_addr_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_addr_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_addr_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_addr_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_addr_s1_readdata),   //                    .readdata
		.out_port   (addr_external_connection_export)       // external_connection.export
	);

	test1a_DONE done (
		.clk      (clk_clk),                            //                 clk.clk
		.reset_n  (~rst_controller_reset_out_reset),    //               reset.reset_n
		.address  (mm_interconnect_0_done_s1_address),  //                  s1.address
		.readdata (mm_interconnect_0_done_s1_readdata), //                    .readdata
		.in_port  (done_external_connection_export)     // external_connection.export
	);

	test1a_ADDR gpio (
		.clk        (clk_clk),                              //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),      //               reset.reset_n
		.address    (mm_interconnect_0_gpio_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_gpio_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_gpio_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_gpio_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_gpio_s1_readdata),   //                    .readdata
		.out_port   (gpio_external_connection_export)       // external_connection.export
	);

	test1a_ADDR led (
		.clk        (clk_clk),                             //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),     //               reset.reset_n
		.address    (mm_interconnect_0_led_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_led_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_led_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_led_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_led_s1_readdata),   //                    .readdata
		.out_port   (led_external_connection_export)       // external_connection.export
	);

	test1a_M_RESET m_reset (
		.clk        (clk_clk),                                 //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),         //               reset.reset_n
		.address    (mm_interconnect_0_m_reset_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_m_reset_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_m_reset_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_m_reset_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_m_reset_s1_readdata),   //                    .readdata
		.out_port   (m_reset_external_connection_export)       // external_connection.export
	);

	test1a_M_RESET oper (
		.clk        (clk_clk),                              //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),      //               reset.reset_n
		.address    (mm_interconnect_0_oper_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_oper_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_oper_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_oper_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_oper_s1_readdata),   //                    .readdata
		.out_port   (oper_external_connection_export)       // external_connection.export
	);

	test1a_M_RESET start (
		.clk        (clk_clk),                               //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),       //               reset.reset_n
		.address    (mm_interconnect_0_start_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_start_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_start_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_start_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_start_s1_readdata),   //                    .readdata
		.out_port   (start_external_connection_export)       // external_connection.export
	);

	test1a_M_RESET start_16 (
		.clk        (clk_clk),                                  //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),          //               reset.reset_n
		.address    (mm_interconnect_0_start_16_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_start_16_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_start_16_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_start_16_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_start_16_s1_readdata),   //                    .readdata
		.out_port   (start_16_external_connection_export)       // external_connection.export
	);

	test1a_WR_DATA wr_data (
		.clk        (clk_clk),                                 //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),         //               reset.reset_n
		.address    (mm_interconnect_0_wr_data_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_wr_data_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_wr_data_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_wr_data_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_wr_data_s1_readdata),   //                    .readdata
		.out_port   (wr_data_external_connection_export)       // external_connection.export
	);

	test1a_WR_DATA_16 wr_data_16 (
		.clk        (clk_clk),                                    //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),            //               reset.reset_n
		.address    (mm_interconnect_0_wr_data_16_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_wr_data_16_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_wr_data_16_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_wr_data_16_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_wr_data_16_s1_readdata),   //                    .readdata
		.out_port   (wr_data_16_external_connection_export)       // external_connection.export
	);

	test1a_master_0 #(
		.USE_PLI     (0),
		.PLI_PORT    (50000),
		.FIFO_DEPTHS (2)
	) master_0 (
		.clk_clk              (clk_clk),                       //          clk.clk
		.clk_reset_reset      (~reset_reset_n),                //    clk_reset.reset
		.master_address       (master_0_master_address),       //       master.address
		.master_readdata      (master_0_master_readdata),      //             .readdata
		.master_read          (master_0_master_read),          //             .read
		.master_write         (master_0_master_write),         //             .write
		.master_writedata     (master_0_master_writedata),     //             .writedata
		.master_waitrequest   (master_0_master_waitrequest),   //             .waitrequest
		.master_readdatavalid (master_0_master_readdatavalid), //             .readdatavalid
		.master_byteenable    (master_0_master_byteenable),    //             .byteenable
		.master_reset_reset   ()                               // master_reset.reset
	);

	test1a_mm_interconnect_0 mm_interconnect_0 (
		.clk_0_clk_clk                                  (clk_clk),                                    //                                clk_0_clk.clk
		.LED_reset_reset_bridge_in_reset_reset          (rst_controller_reset_out_reset),             //          LED_reset_reset_bridge_in_reset.reset
		.master_0_clk_reset_reset_bridge_in_reset_reset (rst_controller_reset_out_reset),             // master_0_clk_reset_reset_bridge_in_reset.reset
		.master_0_master_address                        (master_0_master_address),                    //                          master_0_master.address
		.master_0_master_waitrequest                    (master_0_master_waitrequest),                //                                         .waitrequest
		.master_0_master_byteenable                     (master_0_master_byteenable),                 //                                         .byteenable
		.master_0_master_read                           (master_0_master_read),                       //                                         .read
		.master_0_master_readdata                       (master_0_master_readdata),                   //                                         .readdata
		.master_0_master_readdatavalid                  (master_0_master_readdatavalid),              //                                         .readdatavalid
		.master_0_master_write                          (master_0_master_write),                      //                                         .write
		.master_0_master_writedata                      (master_0_master_writedata),                  //                                         .writedata
		.ADDR_s1_address                                (mm_interconnect_0_addr_s1_address),          //                                  ADDR_s1.address
		.ADDR_s1_write                                  (mm_interconnect_0_addr_s1_write),            //                                         .write
		.ADDR_s1_readdata                               (mm_interconnect_0_addr_s1_readdata),         //                                         .readdata
		.ADDR_s1_writedata                              (mm_interconnect_0_addr_s1_writedata),        //                                         .writedata
		.ADDR_s1_chipselect                             (mm_interconnect_0_addr_s1_chipselect),       //                                         .chipselect
		.DONE_s1_address                                (mm_interconnect_0_done_s1_address),          //                                  DONE_s1.address
		.DONE_s1_readdata                               (mm_interconnect_0_done_s1_readdata),         //                                         .readdata
		.GPIO_s1_address                                (mm_interconnect_0_gpio_s1_address),          //                                  GPIO_s1.address
		.GPIO_s1_write                                  (mm_interconnect_0_gpio_s1_write),            //                                         .write
		.GPIO_s1_readdata                               (mm_interconnect_0_gpio_s1_readdata),         //                                         .readdata
		.GPIO_s1_writedata                              (mm_interconnect_0_gpio_s1_writedata),        //                                         .writedata
		.GPIO_s1_chipselect                             (mm_interconnect_0_gpio_s1_chipselect),       //                                         .chipselect
		.LED_s1_address                                 (mm_interconnect_0_led_s1_address),           //                                   LED_s1.address
		.LED_s1_write                                   (mm_interconnect_0_led_s1_write),             //                                         .write
		.LED_s1_readdata                                (mm_interconnect_0_led_s1_readdata),          //                                         .readdata
		.LED_s1_writedata                               (mm_interconnect_0_led_s1_writedata),         //                                         .writedata
		.LED_s1_chipselect                              (mm_interconnect_0_led_s1_chipselect),        //                                         .chipselect
		.M_RESET_s1_address                             (mm_interconnect_0_m_reset_s1_address),       //                               M_RESET_s1.address
		.M_RESET_s1_write                               (mm_interconnect_0_m_reset_s1_write),         //                                         .write
		.M_RESET_s1_readdata                            (mm_interconnect_0_m_reset_s1_readdata),      //                                         .readdata
		.M_RESET_s1_writedata                           (mm_interconnect_0_m_reset_s1_writedata),     //                                         .writedata
		.M_RESET_s1_chipselect                          (mm_interconnect_0_m_reset_s1_chipselect),    //                                         .chipselect
		.OPER_s1_address                                (mm_interconnect_0_oper_s1_address),          //                                  OPER_s1.address
		.OPER_s1_write                                  (mm_interconnect_0_oper_s1_write),            //                                         .write
		.OPER_s1_readdata                               (mm_interconnect_0_oper_s1_readdata),         //                                         .readdata
		.OPER_s1_writedata                              (mm_interconnect_0_oper_s1_writedata),        //                                         .writedata
		.OPER_s1_chipselect                             (mm_interconnect_0_oper_s1_chipselect),       //                                         .chipselect
		.START_s1_address                               (mm_interconnect_0_start_s1_address),         //                                 START_s1.address
		.START_s1_write                                 (mm_interconnect_0_start_s1_write),           //                                         .write
		.START_s1_readdata                              (mm_interconnect_0_start_s1_readdata),        //                                         .readdata
		.START_s1_writedata                             (mm_interconnect_0_start_s1_writedata),       //                                         .writedata
		.START_s1_chipselect                            (mm_interconnect_0_start_s1_chipselect),      //                                         .chipselect
		.START_16_s1_address                            (mm_interconnect_0_start_16_s1_address),      //                              START_16_s1.address
		.START_16_s1_write                              (mm_interconnect_0_start_16_s1_write),        //                                         .write
		.START_16_s1_readdata                           (mm_interconnect_0_start_16_s1_readdata),     //                                         .readdata
		.START_16_s1_writedata                          (mm_interconnect_0_start_16_s1_writedata),    //                                         .writedata
		.START_16_s1_chipselect                         (mm_interconnect_0_start_16_s1_chipselect),   //                                         .chipselect
		.WR_DATA_s1_address                             (mm_interconnect_0_wr_data_s1_address),       //                               WR_DATA_s1.address
		.WR_DATA_s1_write                               (mm_interconnect_0_wr_data_s1_write),         //                                         .write
		.WR_DATA_s1_readdata                            (mm_interconnect_0_wr_data_s1_readdata),      //                                         .readdata
		.WR_DATA_s1_writedata                           (mm_interconnect_0_wr_data_s1_writedata),     //                                         .writedata
		.WR_DATA_s1_chipselect                          (mm_interconnect_0_wr_data_s1_chipselect),    //                                         .chipselect
		.WR_DATA_16_s1_address                          (mm_interconnect_0_wr_data_16_s1_address),    //                            WR_DATA_16_s1.address
		.WR_DATA_16_s1_write                            (mm_interconnect_0_wr_data_16_s1_write),      //                                         .write
		.WR_DATA_16_s1_readdata                         (mm_interconnect_0_wr_data_16_s1_readdata),   //                                         .readdata
		.WR_DATA_16_s1_writedata                        (mm_interconnect_0_wr_data_16_s1_writedata),  //                                         .writedata
		.WR_DATA_16_s1_chipselect                       (mm_interconnect_0_wr_data_16_s1_chipselect)  //                                         .chipselect
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller (
		.reset_in0      (~reset_reset_n),                 // reset_in0.reset
		.clk            (clk_clk),                        //       clk.clk
		.reset_out      (rst_controller_reset_out_reset), // reset_out.reset
		.reset_req      (),                               // (terminated)
		.reset_req_in0  (1'b0),                           // (terminated)
		.reset_in1      (1'b0),                           // (terminated)
		.reset_req_in1  (1'b0),                           // (terminated)
		.reset_in2      (1'b0),                           // (terminated)
		.reset_req_in2  (1'b0),                           // (terminated)
		.reset_in3      (1'b0),                           // (terminated)
		.reset_req_in3  (1'b0),                           // (terminated)
		.reset_in4      (1'b0),                           // (terminated)
		.reset_req_in4  (1'b0),                           // (terminated)
		.reset_in5      (1'b0),                           // (terminated)
		.reset_req_in5  (1'b0),                           // (terminated)
		.reset_in6      (1'b0),                           // (terminated)
		.reset_req_in6  (1'b0),                           // (terminated)
		.reset_in7      (1'b0),                           // (terminated)
		.reset_req_in7  (1'b0),                           // (terminated)
		.reset_in8      (1'b0),                           // (terminated)
		.reset_req_in8  (1'b0),                           // (terminated)
		.reset_in9      (1'b0),                           // (terminated)
		.reset_req_in9  (1'b0),                           // (terminated)
		.reset_in10     (1'b0),                           // (terminated)
		.reset_req_in10 (1'b0),                           // (terminated)
		.reset_in11     (1'b0),                           // (terminated)
		.reset_req_in11 (1'b0),                           // (terminated)
		.reset_in12     (1'b0),                           // (terminated)
		.reset_req_in12 (1'b0),                           // (terminated)
		.reset_in13     (1'b0),                           // (terminated)
		.reset_req_in13 (1'b0),                           // (terminated)
		.reset_in14     (1'b0),                           // (terminated)
		.reset_req_in14 (1'b0),                           // (terminated)
		.reset_in15     (1'b0),                           // (terminated)
		.reset_req_in15 (1'b0)                            // (terminated)
	);

endmodule
